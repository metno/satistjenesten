netcdf amsr2n90 {
dimensions:
	time = 1 ;
	ni = 5 ;
	nih = 5 ;
	n85 = 4 ;
variables:
	double time(time) ;
		time:_FillValue = -10000000000. ;
		time:units = "seconds since 2010-01-01 00:00:00" ;
		time:long_name = "reference time of swath data" ;
	float lat_l(ni) ;
		lat_l:_FillValue = -1.e+10f ;
		lat_l:units = "degrees_north" ;
		lat_l:long_name = "latitude low res obs" ;
	float lon_l(ni) ;
		lon_l:_FillValue = -1.e+10f ;
		lon_l:units = "degrees_east" ;
		lon_l:long_name = "longitude low res obs" ;
	short dtime(ni) ;
		dtime:_FillValue = -32767s ;
		dtime:units = "second" ;
		dtime:long_name = "time difference from reference time" ;
		dtime:scale_factor = 1.f ;
	short surf_l(ni) ;
		surf_l:_FillValue = -32767s ;
		surf_l:units = "1" ;
		surf_l:long_name = "surface flag, low res obs" ;
		surf_l:coordinates = "dtime lat_l lon_l" ;
		surf_l:comment = "-1 = unknown, 0 = land, 2 = near coast, 3 = ice shelves/land ice, 4 = possible ice, 5 = ice-free ocean, 6 = coast" ;
	float tb19v(ni) ;
		tb19v:_FillValue = -1.e+10f ;
		tb19v:units = "K" ;
		tb19v:long_name = "BT 19V GHz" ;
		tb19v:coordinates = "dtime lat_l lon_l" ;
	float tb19h(ni) ;
		tb19h:_FillValue = -1.e+10f ;
		tb19h:units = "K" ;
		tb19h:long_name = "BT 19H GHz" ;
	float tb37v(ni) ;
		tb37v:_FillValue = -1.e+10f ;
		tb37v:units = "K" ;
		tb37v:long_name = "BT 37V GHz" ;
		tb37v:coordinates = "dtime lat_l lon_l" ;
	float tb37h(ni) ;
		tb37h:_FillValue = -1.e+10f ;
		tb37h:units = "K" ;
		tb37h:long_name = "BT 37H GHz" ;
	float tb22(ni) ;
		tb22:_FillValue = -1.e+10f ;
		tb22:units = "K" ;
		tb22:long_name = "BT 22V GHz" ;
		tb22:coordinates = "dtime lat_l lon_l" ;
	float lat_h(nih, n85) ;
		lat_h:_FillValue = -1.e+10f ;
		lat_h:units = "degrees_north" ;
		lat_h:long_name = "latitude high res obs" ;
	float lon_h(nih, n85) ;
		lon_h:_FillValue = -1.e+10f ;
		lon_h:units = "degrees_east" ;
		lon_h:long_name = "longitude high res obs" ;
	short surf_h(nih, n85) ;
		surf_h:_FillValue = -32767s ;
		surf_h:units = "1" ;
		surf_h:long_name = "surface flag, high res obs" ;
		surf_h:coordinates = "dtime_h lat_h lon_h" ;
	float tb85v(nih, n85) ;
		tb85v:_FillValue = -1.e+10f ;
		tb85v:units = "K" ;
		tb85v:long_name = "BT 85V GHz" ;
		tb85v:coordinates = "dtime_h lat_h lon_h" ;
	float tb85h(nih, n85) ;
		tb85h:_FillValue = -1.e+10f ;
		tb85h:units = "K" ;
		tb85h:long_name = "BT 85H GHz" ;
		tb85h:coordinates = "dtime_h lat_h lon_h" ;
	short ct_NASA(ni) ;
		ct_NASA:_FillValue = -32767s ;
		ct_NASA:units = "%" ;
		ct_NASA:long_name = "Uncorrected total ice concentration using NASA Team" ;
		ct_NASA:scale_factor = 0.01f ;
	byte wf_NASA(ni) ;
		wf_NASA:_FillValue = -1b ;
		wf_NASA:units = "1" ;
		wf_NASA:long_name = "Weather filter from Cavalieri et al. (1992)" ;
		wf_NASA:comment = "1: Probably OW, 0: Probably ICE" ;
	short ct_NASA_wWF(ni) ;
		ct_NASA_wWF:_FillValue = -32767s ;
		ct_NASA_wWF:units = "%" ;
		ct_NASA_wWF:long_name = "Uncorrected total ice concentration using NASA Team, screened by Weather Filter" ;
		ct_NASA_wWF:scale_factor = 0.01f ;
	short wind_speed(ni) ;
		wind_speed:_FillValue = -32767s ;
		wind_speed:units = "m/s" ;
		wind_speed:long_name = "NWP 10m wind speed" ;
		wind_speed:scale_factor = 0.01f ;
	short air_temp(ni) ;
		air_temp:_FillValue = -32767s ;
		air_temp:units = "K" ;
		air_temp:long_name = "NWP air temperature (at 2m)" ;
		air_temp:scale_factor = 0.01f ;
		air_temp:add_offset = 273 ;
	short tcwv(ni) ;
		tcwv:_FillValue = -32767s ;
		tcwv:units = "kg/m2" ;
		tcwv:long_name = "NWP total column water vapour" ;
		tcwv:scale_factor = 0.01f ;
	short dtb19v_OSISAF_corrNASA(ni) ;
		dtb19v_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb19v_OSISAF_corrNASA:units = "K" ;
		dtb19v_OSISAF_corrNASA:long_name = "correction of BT 19v GHz using NASA Team" ;
		dtb19v_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb19h_OSISAF_corrNASA(ni) ;
		dtb19h_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb19h_OSISAF_corrNASA:units = "K" ;
		dtb19h_OSISAF_corrNASA:long_name = "correction of BT 19h GHz using NASA Team" ;
		dtb19h_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb22v_OSISAF_corrNASA(ni) ;
		dtb22v_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb22v_OSISAF_corrNASA:units = "K" ;
		dtb22v_OSISAF_corrNASA:long_name = "correction of BT 22v GHz using NASA Team" ;
		dtb22v_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb22h_OSISAF_corrNASA(ni) ;
		dtb22h_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb22h_OSISAF_corrNASA:units = "K" ;
		dtb22h_OSISAF_corrNASA:long_name = "correction of BT 22h GHz using NASA Team" ;
		dtb22h_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb37v_OSISAF_corrNASA(ni) ;
		dtb37v_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb37v_OSISAF_corrNASA:units = "K" ;
		dtb37v_OSISAF_corrNASA:long_name = "correction of BT 37v GHz using NASA Team" ;
		dtb37v_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb37h_OSISAF_corrNASA(ni) ;
		dtb37h_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb37h_OSISAF_corrNASA:units = "K" ;
		dtb37h_OSISAF_corrNASA:long_name = "correction of BT 37h GHz using NASA Team" ;
		dtb37h_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb85h_OSISAF_corrNASA(ni, n85) ;
		dtb85h_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb85h_OSISAF_corrNASA:units = "K" ;
		dtb85h_OSISAF_corrNASA:long_name = "correction of BT 85h GHz using NASA Team" ;
		dtb85h_OSISAF_corrNASA:scale_factor = 0.01f ;
	short dtb85v_OSISAF_corrNASA(ni, n85) ;
		dtb85v_OSISAF_corrNASA:_FillValue = -32767s ;
		dtb85v_OSISAF_corrNASA:units = "K" ;
		dtb85v_OSISAF_corrNASA:long_name = "correction of BT 85v GHz using NASA Team" ;
		dtb85v_OSISAF_corrNASA:scale_factor = 0.01f ;
	short ct_OSISAF_corrNASA(ni) ;
		ct_OSISAF_corrNASA:_FillValue = -32767s ;
		ct_OSISAF_corrNASA:units = "%" ;
		ct_OSISAF_corrNASA:long_name = "OSISAF ice concentration using NASA brightness temperatures and tie-points" ;
		ct_OSISAF_corrNASA:scale_factor = 0.01f ;
	short ct_n90_OSISAF_corrNASA(ni, n85) ;
		ct_n90_OSISAF_corrNASA:_FillValue = -32767s ;
		ct_n90_OSISAF_corrNASA:units = "%" ;
		ct_n90_OSISAF_corrNASA:long_name = "OSISAF n90 ice concentration using NASA brightness temperatures and tie-points" ;
		ct_n90_OSISAF_corrNASA:scale_factor = 0.01f ;
	byte wf_NASA_n90(ni, n85) ;
		wf_NASA_n90:_FillValue = -1b ;
	short ct_n90_OSISAF_corrNASA_wWF(ni, n85) ;
		ct_n90_OSISAF_corrNASA_wWF:_FillValue = -32767s ;
		ct_n90_OSISAF_corrNASA_wWF:units = "%" ;
		ct_n90_OSISAF_corrNASA_wWF:long_name = "OSISAF ice concentration using NASA brightness temperatures and tie-points, screened by Weather Filter" ;
		ct_n90_OSISAF_corrNASA_wWF:scale_factor = 0.01f ;

// global attributes:
		:title = "L1 amsr satellite data" ;
		:Conventions = "CF-1.0" ;
		:institution = "Ocean and Sea Ice Satellite Application Facility (OSI SAF)" ;
		:orbit_number = -999. ;
		:satellite = "gw1" ;
		:start_date_and_time = "2015-03-30T10:04:04Z" ;
		:end_date_and_time = "2015-03-30T11:40:02Z" ;
		:history = "Created 2015-03-30" ;
		:fromfile = "GW1AM2_201503301003_046B_L1SNBTBR_2200200.h5" ;
		:scanline_length = 243 ;
}
